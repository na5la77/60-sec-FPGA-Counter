version https://git-lfs.github.com/spec/v1
oid sha256:46a7cdf5fe8a14738cf2fa3a60335a04f1d7a85af193cfdb5e8932a5cd76b2d6
size 831
