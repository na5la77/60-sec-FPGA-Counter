version https://git-lfs.github.com/spec/v1
oid sha256:4fe3e8d0ed8fb16bb2bdeb85efd58c3a5b0a2167a8c4669be59dd29fbc53511e
size 3659
