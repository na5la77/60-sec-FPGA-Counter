version https://git-lfs.github.com/spec/v1
oid sha256:ce7496dd90eb36b547b3e2c8d05c0bc173dc0c55d960c49128cd774fe86ee43d
size 726
