version https://git-lfs.github.com/spec/v1
oid sha256:b08478d5513d57dbf267e3394d5b30b572c486f88a342b740f750f9dad65e2c9
size 751
