version https://git-lfs.github.com/spec/v1
oid sha256:e5d2a553988de2df682c6d676fd0e4c7f8ac5ba958204d4f0e3292c52f10b0f7
size 775
