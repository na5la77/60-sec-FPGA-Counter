version https://git-lfs.github.com/spec/v1
oid sha256:b08ef553ad5a2bd0bce29078105b5d728feec4c353f4a84fad64b743c7902a65
size 1074
